module sjosj 12311