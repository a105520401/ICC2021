module sjosj